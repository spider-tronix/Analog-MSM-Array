magic
tech sky130A
timestamp 1646067201
<< nmos >>
rect 0 0 15 2500
rect 145 0 160 2500
rect 290 0 305 2500
rect 435 0 450 2500
rect 580 0 595 2500
rect 725 0 740 2500
rect 870 0 885 2500
rect 1015 0 1030 2500
rect 1160 0 1175 2500
rect 1305 0 1320 2500
<< ndiff >>
rect -50 2485 0 2500
rect -50 15 -35 2485
rect -15 15 0 2485
rect -50 0 0 15
rect 15 2485 65 2500
rect 15 15 30 2485
rect 50 15 65 2485
rect 15 0 65 15
rect 95 2485 145 2500
rect 95 15 110 2485
rect 130 15 145 2485
rect 95 0 145 15
rect 160 2485 210 2500
rect 160 15 175 2485
rect 195 15 210 2485
rect 160 0 210 15
rect 240 2485 290 2500
rect 240 15 255 2485
rect 275 15 290 2485
rect 240 0 290 15
rect 305 2485 355 2500
rect 305 15 320 2485
rect 340 15 355 2485
rect 305 0 355 15
rect 385 2485 435 2500
rect 385 15 400 2485
rect 420 15 435 2485
rect 385 0 435 15
rect 450 2485 500 2500
rect 450 15 465 2485
rect 485 15 500 2485
rect 450 0 500 15
rect 530 2485 580 2500
rect 530 15 545 2485
rect 565 15 580 2485
rect 530 0 580 15
rect 595 2485 645 2500
rect 595 15 610 2485
rect 630 15 645 2485
rect 595 0 645 15
rect 675 2485 725 2500
rect 675 15 690 2485
rect 710 15 725 2485
rect 675 0 725 15
rect 740 2485 790 2500
rect 740 15 755 2485
rect 775 15 790 2485
rect 740 0 790 15
rect 820 2485 870 2500
rect 820 15 835 2485
rect 855 15 870 2485
rect 820 0 870 15
rect 885 2485 935 2500
rect 885 15 900 2485
rect 920 15 935 2485
rect 885 0 935 15
rect 965 2485 1015 2500
rect 965 15 980 2485
rect 1000 15 1015 2485
rect 965 0 1015 15
rect 1030 2485 1080 2500
rect 1030 15 1045 2485
rect 1065 15 1080 2485
rect 1030 0 1080 15
rect 1110 2485 1160 2500
rect 1110 15 1125 2485
rect 1145 15 1160 2485
rect 1110 0 1160 15
rect 1175 2485 1225 2500
rect 1175 15 1190 2485
rect 1210 15 1225 2485
rect 1175 0 1225 15
rect 1255 2485 1305 2500
rect 1255 15 1270 2485
rect 1290 15 1305 2485
rect 1255 0 1305 15
rect 1320 2485 1370 2500
rect 1320 15 1335 2485
rect 1355 15 1370 2485
rect 1320 0 1370 15
<< ndiffc >>
rect -35 15 -15 2485
rect 30 15 50 2485
rect 110 15 130 2485
rect 175 15 195 2485
rect 255 15 275 2485
rect 320 15 340 2485
rect 400 15 420 2485
rect 465 15 485 2485
rect 545 15 565 2485
rect 610 15 630 2485
rect 690 15 710 2485
rect 755 15 775 2485
rect 835 15 855 2485
rect 900 15 920 2485
rect 980 15 1000 2485
rect 1045 15 1065 2485
rect 1125 15 1145 2485
rect 1190 15 1210 2485
rect 1270 15 1290 2485
rect 1335 15 1355 2485
<< psubdiff >>
rect -100 2485 -50 2500
rect -100 15 -85 2485
rect -65 15 -50 2485
rect -100 0 -50 15
<< psubdiffcont >>
rect -85 15 -65 2485
<< poly >>
rect 0 2500 15 2515
rect 145 2500 160 2515
rect 290 2500 305 2515
rect 435 2500 450 2515
rect 580 2500 595 2515
rect 725 2500 740 2515
rect 870 2500 885 2515
rect 1015 2500 1030 2515
rect 1160 2500 1175 2515
rect 1305 2500 1320 2515
rect 0 -15 15 0
rect 145 -15 160 0
rect 290 -15 305 0
rect 435 -15 450 0
rect 580 -15 595 0
rect 725 -15 740 0
rect 870 -15 885 0
rect 1015 -15 1030 0
rect 1160 -15 1175 0
rect 1305 -15 1320 0
<< locali >>
rect -95 2485 -5 2495
rect -95 15 -85 2485
rect -65 15 -35 2485
rect -15 15 -5 2485
rect -95 5 -5 15
rect 20 2485 60 2495
rect 20 15 30 2485
rect 50 15 60 2485
rect 20 5 60 15
rect 95 2485 140 2495
rect 95 15 110 2485
rect 130 15 140 2485
rect 95 5 140 15
rect 165 2485 205 2495
rect 165 15 175 2485
rect 195 15 205 2485
rect 165 5 205 15
rect 240 2485 285 2495
rect 240 15 255 2485
rect 275 15 285 2485
rect 240 5 285 15
rect 310 2485 350 2495
rect 310 15 320 2485
rect 340 15 350 2485
rect 310 5 350 15
rect 385 2485 430 2495
rect 385 15 400 2485
rect 420 15 430 2485
rect 385 5 430 15
rect 455 2485 495 2495
rect 455 15 465 2485
rect 485 15 495 2485
rect 455 5 495 15
rect 530 2485 575 2495
rect 530 15 545 2485
rect 565 15 575 2485
rect 530 5 575 15
rect 600 2485 640 2495
rect 600 15 610 2485
rect 630 15 640 2485
rect 600 5 640 15
rect 675 2485 720 2495
rect 675 15 690 2485
rect 710 15 720 2485
rect 675 5 720 15
rect 745 2485 785 2495
rect 745 15 755 2485
rect 775 15 785 2485
rect 745 5 785 15
rect 820 2485 865 2495
rect 820 15 835 2485
rect 855 15 865 2485
rect 820 5 865 15
rect 890 2485 930 2495
rect 890 15 900 2485
rect 920 15 930 2485
rect 890 5 930 15
rect 965 2485 1010 2495
rect 965 15 980 2485
rect 1000 15 1010 2485
rect 965 5 1010 15
rect 1035 2485 1075 2495
rect 1035 15 1045 2485
rect 1065 15 1075 2485
rect 1035 5 1075 15
rect 1110 2485 1155 2495
rect 1110 15 1125 2485
rect 1145 15 1155 2485
rect 1110 5 1155 15
rect 1180 2485 1220 2495
rect 1180 15 1190 2485
rect 1210 15 1220 2485
rect 1180 5 1220 15
rect 1255 2485 1300 2495
rect 1255 15 1270 2485
rect 1290 15 1300 2485
rect 1255 5 1300 15
rect 1325 2485 1365 2495
rect 1325 15 1335 2485
rect 1355 15 1365 2485
rect 1325 5 1365 15
<< end >>
